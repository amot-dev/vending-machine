ENTITY programmingUnit IS
PORT (clock, reset, hardReset, set, enable : IN STD_LOGIC;
		product										 : IN UNSIGNED(1 DOWNTO 0);
		QDN											 : IN STD_LOGic_VECTOR(2 DOWNTO 0);
		writeEnable									 : OUT STD_LOGIC;
		data, address								 : OUT UNSIGNED(5 DOWNTO 0));
END programmingUnit;

ARCHITECTURE Behaviour OF programmingUnit IS

BEGIN
END Behaviour;
